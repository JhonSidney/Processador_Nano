module 

endmodule 