module
endmodule 